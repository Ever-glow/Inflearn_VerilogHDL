//////////////////////////////////////////////////////////////////////////////////
// Company: Personal
// Engineer: Matbi / Austin
//
// Create Date:
// Design Name: hello_world
// Module Name: hello_world
// Project Name:
// Target Devices:
// Tool Versions:
// Description: hello_world test
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module hello_world;

initial begin
$display("hello world");
$finish;
end

endmodule
